//`timescale 1ns / 1ps

//module movement(
//	input CLK100MHZ,
//    input reset,
//    input [2:0] movementCommand, 
//    input [1:0] speed,
//    input [1:0] speedChange,
//    output enableA,
//    output enableB,
//    output [3:0] motor
//    );
//    always @(*) begin 
//    //foo
//    end
//endmodule
