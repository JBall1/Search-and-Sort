`timescale 1ns / 1ps

module metalDetector(
        input CLK100MHZ
        //input metalVal,
        //output metalFlagt
    );
    
    
always @ (posedge CLK100MHZ) begin
       
//       if (metalVal < 1) begin
//         metalFlagt = 0;
//       end
       
//       else if (metalVal >= 1) begin
//         metalFlagt <= 1;
//       end
       
//       end
end
endmodule
